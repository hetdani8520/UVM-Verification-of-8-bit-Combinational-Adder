`include "comb_adder_item.sv"
`include "agent_config.sv"
`include "env_config.sv"
`include "comb_adder_seq.sv"
`include "adder_driver.sv"
`include "adder_monitor.sv"
`include "adder_scb.sv"
`include "adder_predictor.sv"
`include "adder_agent.sv"
`include "adder_env.sv"